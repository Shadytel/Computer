----------------------------------------------------------------------------------
-- Company: Lake Union Bell
-- Engineer: Nick Burrows
-- 
-- Create Date:    19:49:20 09/22/2011 
-- Design Name: 
-- Module Name:    RAM - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

library UNISIM;
use UNISIM.VComponents.all;

entity RAM is
  Port
		(
			CLK: in std_logic;
			Control: in std_logic_vector(11 downto 0);
			ADDR: in std_logic_vector(11 downto 0);
			IO: inout std_logic_vector(11 downto 0)
		);

end RAM;

architecture Behavioral of RAM is
 signal SSR: std_logic; 
 signal RAMBus: std_logic_vector(11 downto 0) := "000000000000";
begin
    SSR <= '0';
	 
	 process (Control, RAMBus)
	 begin
		if(Control(0) = '1') then
			IO <= RAMBus;
		else
			IO <= "ZZZZZZZZZZZZ";
		end if;
	 end process;
	
	 
	 LowNibble : RAMB16_S4 
		generic map ( 
				INIT => X"A", --  Value of output RAM registers at startup
				SRVAL => X"0", --  Ouput value upon SSR assertion
				WRITE_MODE => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
				INIT_00 => X"F00000000000000000000000000000000000A010F5E460F00000000051100001", --Ram contents in hex, higher addresses right most
				INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
				-- Address 1024 to 2047
				INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
				-- Address 2048 to 3071
				INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
				-- Address 3072 to 4095
				INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")							
			port map (
				DO => RAMBus(3 downto 0),      -- 4-bit Data Output
				ADDR =>  ADDR,  -- 12-bit Address Input
				CLK => CLK,    -- Clock
				DI => IO(3 downto 0),      -- 4-bit Data Input
				EN => '1',      -- RAM Enable Input
				SSR => SSR,    -- Synchronous Set/Reset Input
				WE => Control(1) -- Write Enable Input
		);
		
	MiddleNibble : RAMB16_S4 
		generic map ( 
				INIT => X"1", --  Value of output RAM registers at startup
				SRVAL => X"0", --  Ouput value upon SSR assertion
				WRITE_MODE => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
				INIT_00 => X"C000000000000000000000000000000000001010F2230CF00000000000000001",
				INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
				-- Address 1024 to 2047
				INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
				-- Address 2048 to 3071
				INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
				-- Address 3072 to 4095
				INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")		
			port map (
				DO => RAMBus(7 downto 4),      -- 4-bit Data Output
				ADDR =>  ADDR,  -- 12-bit Address Input
				CLK => CLK,    -- Clock
				DI => IO(7 downto 4),      -- 4-bit Data Input
				EN => '1',      -- RAM Enable Input
				SSR => SSR,    -- Synchronous Set/Reset Input
				WE => Control(1)       -- Write Enable Input
		);
		
	HighNibble : RAMB16_S4 
		generic map ( 
				INIT => X"0", --  Value of output RAM registers at startup
				SRVAL => X"0", --  Ouput value upon SSR assertion
				WRITE_MODE => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
				INIT_00 => X"D000000000000000000000000000000000000A0A08080D700000000000000000",
				INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
				-- Address 1024 to 2047
				INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
				-- Address 2048 to 3071
				INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
				-- Address 3072 to 4095
				INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")				
			port map (
				DO => RAMBus(11 downto 8),      -- 4-bit Data Output
				ADDR =>  ADDR,  -- 12-bit Address Input
				CLK => CLK,    -- Clock
				DI => IO(11 downto 8),      -- 4-bit Data Input
				EN => '1',      -- RAM Enable Input
				SSR => SSR,    -- Synchronous Set/Reset Input
				WE => Control(1)      -- Write Enable Input
		);
  
  
end Behavioral;

